package lc3_prediction_pkg;
   import uvm_pkg::*;

   `include "src/lc3_prediction_typedefs.svh"
   `include "src/fetch_model.svh"
   `include "src/decode_model.svh"
   `include "src/execute_model.svh"
   `include "src/mem_access_model.svh"
   `include "src/writeback_model.svh"
   `include "src/controller_model.svh"

endpackage
